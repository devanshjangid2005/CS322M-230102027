module Q2(
    input [3:0] A,
    input [3:0] B,
    output C
);

assign C=(A==B);

endmodule
